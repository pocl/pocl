package tta_core_imem_mau is
   -- created by generatebits
   constant IMEMMAUWIDTH : positive := 42;
end tta_core_imem_mau;

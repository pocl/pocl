library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use work.tta_core_imem_mau.all;

package tta_core_imem_image is

  type std_logic_imem_matrix is array (natural range <>) of std_logic_vector(IMEMMAUWIDTH-1 downto 0);

  constant imem_array : std_logic_imem_matrix := (
"000000000000000000000000000000000100111000",
"000110000000000000000000000000000000111100",
"000000000000000000000000000000000110110010",
"000000000000000000000000001110000000001000",
"000101100000000000000000000000000000010000",
"000101100000000000000000000000000000101110",
"000000000000000000000000000000000000010101",
"000000000000000000000000000000000100111000",
"000100000000000000000000000000000000001000",
"000110000000000000000000000000000000111100",
"000101100000000000000000000000000000101110",
"000000000000000000000000000001011000111000",
"000101100000000000000000000000000000001000",
"000101100000000000000000000000000000010000",
"000101100000000000000000000000000000111000",
"000000000000000000000000000000100101110011",
"000000000000000000000000000001010100000000",
"000100000000000000000000000000000010111100",
"000101100000000000000000000000000000101110",
"000100000000000000000000000000000000111000",
"000000000000000000000000000000001100000000",
"000101100000000000000000000000000000101001",
"101111111111111111111111111111111111111111",
"000000000000000000000000000000000001110101",
"000111000000000000000000000000000000111000",
"000000000000000000000000000000111000000000",
"000101100000000000000000000000000000101001",
"000000000000000000000000000000000001111100",
"000111000000000000000000000000000000101101",
"000100000000000000000000000000000000111000",
"000000000000000000000000000000001000000000",
"000101100000000000000000000000000000101001",
"000000000000000000000000000000000001110110",
"000111000000000000000000000000000000100110",
"000111000000000000000000000000000000111000",
"000000000000000000000000000000000001000000",
"000101100000000000000000000000000000010101",
"000100000000000000000000000000000000111000",
"000000000000000000000000000000001000000000",
"000100000000000000000000000000000101111100",
"000101100000000000000000000000000000101110",
"000100000000000000000000000000000101111000",
"000100000000000000000000000000000101000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000000000000000000000000000001000000000001",
"000101100000000000000000000000000000111000",
"000000000000000000000000001110000000000101",
"000101100000000000000000000000000000011010",
"000100000000000000000000000000001010101011",
"101111111111111111111111111111111111111111",
"101111111111111111111111111111111111111111",
"000111000000000000000000000000000000111000",
"000000000000000000000000000000000001000010",
"000101100000000000000000000000000000110000",
"001000000000000000000000000000111101110011",
"001100000000000000000000000000001010101011",
"101111111111111111111111111111111111111111",
"101111111111111111111111111111111111111111",
"000100000000000000000000000000001010111000",
"000000000000000000000000000000101000000000",
"000101100000000000000000000000000000101001",
"101111111111111111111111111111111111111111",
"101111111111111111111111111111111111111111",
"000111000000000000000000000000000000010111",
"000111000000000000000000000000000000111000",
"000000000000000000000000000000001001000000",
"000101100000000000000000000000000000100100",
"000000000000000000000000000000001000000000",
"000101100000000000000000000000000000100100",
"000101000000000000000000000000000000111000",
"000101000000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101000000000000000000000000000000111000",
"000101100000000000000000000000000000000101",
"000101100000000000000000000000000000010100",
"000111000000000000000000000000000000111000",
"000000000000000000000000000000000101000000",
"000101100000000000000000000000000000100100",
"000000000000000000000000000000000100000000",
"000101100000000000000000000000000000100100",
"000101000000000000000000000000000000111000",
"000101000000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101000000000000000000000000000000111000",
"000101100000000000000000000000000000000101",
"000101100000000000000000000000000000010101",
"000100000000000000000000000000000111111000",
"000000000000000000000000000000000001000000",
"000101100000000000000000000000000000100100",
"101111111111111111111111111111111111111111",
"000100000000000000000000000000000111100100",
"000101000000000000000000000000000000111000",
"000101000000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101000000000000000000000000000000111000",
"000101100000000000000000000000000000000101",
"000101100000000000000000000000000000010110",
"000100000000000000000000000000000111111000",
"000000000000000000000000000000000011000000",
"000101100000000000000000000000000000100010",
"000100000000000000000000000000001010011110",
"000000000000000000000000000000000111000000",
"000101100000000000000000000000000000100010",
"000101000000000000000000000000000000011001",
"000000000000000000000000000000001011000000",
"000101100000000000000000000000000000100010",
"000101000000000000000000000000000000011011",
"000000000000000000000000000000000010000000",
"000101100000000000000000000000000000100100",
"000101000000000000000000000000000000011101",
"000000000000000000000000000000000110000000",
"000101000000000000000000000000000000011100",
"000101100000000000000000000000000000100100",
"000000000000000000000000000000001010000000",
"000101100000000000000000000000000000010111",
"000100000000000000000000000000001010111000",
"000101000000000000000000000000000000011010",
"000000000000000000000000000000001100000000",
"000101100000000000000000000000000000101001",
"000100000000000000000000000000000000111000",
"000000000000000000000000000000010100000000",
"000111000000000000000000000000000000111100",
"000101100000000000000000000000000000101110",
"000000000000000000000000000000001100000000",
"000101100000000000000000000000000000010010",
"000100000000000000000000000000000111100100",
"000100000000000000000000000000001110111100",
"000100000000000000000000000000001110111000",
"000000000000000000000000000000000010000000",
"000101100000000000000000000000000000101011",
"000101100000000000000000000000000000010111",
"000100000000000000000000000000000010101110",
"000111000000000000000000000000000000111000",
"000000000000000000000000000000000010000100",
"000101100000000000000000000000000000110000",
"000101000000000000000000000000000000111000",
"000101000000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000011000",
"000100000000000000000000000000001100111000",
"000100000000000000000000000000001100000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000011100",
"000100000000000000000000000000001010111000",
"000100000000000000000000000000001010000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000011010",
"000100000000000000000000000000001001111000",
"000100000000000000000000000000001001000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000011110",
"000100000000000000000000000000000000111000",
"000000000000000000000000000000110100000000",
"000000000000000000000000000000000001111100",
"000101100000000000000000000000000000101110",
"000100000000000000000000000000001011111000",
"000100000000000000000000000000001011000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000011011",
"000100000000000000000000000000001101111000",
"000100000000000000000000000000001101000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"001000000000000000000000000110111001110011",
"000101100000000000000000000000000000111000",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000011101",
"000100000000000000000000000000000000111000",
"000000000000000000000000000000001100000000",
"000101100000000000000000000000000000101001",
"101111111111111111111111111111111111111111",
"101111111111111111111111111111111111111111",
"000111000000000000000000000000000000111000",
"000000000000000000000000000000010000000000",
"000101100000000000000000000000000000101001",
"000100000000000000000000000000000000111000",
"000000000000000000000000000000110100000000",
"000111000000000000000000000000000000111100",
"000101100000000000000000000000000000101110",
"000100000000000000000000000000000000111000",
"000000000000000000000000000000110000000000",
"000101100000000000000000000000000000010010",
"000100000000000000000000000000001010111000",
"000100000000000000000000000000000101000101",
"000101100000000000000000000000000000010101",
"000100000000000000000000000000001110111000",
"000100000000000000000000000000001110000000",
"000101100000000000000000000000000000011010",
"000100000000000000000000000000001011111000",
"000100000000000000000000000000001011000000",
"000101100000000000000000000000000000011001",
"000100000000000000000000000000001000111000",
"000100000000000000000000000000000100000101",
"000101100000000000000000000000000000010100",
"000100000000000000000000000000001101111000",
"000100000000000000000000000000001101000000",
"000101100000000000000000000000000000011000",
"000100000000000000000000000000001100111000",
"000100000000000000000000000000000110000101",
"000100000000000000000000000000000111101011",
"000101100000000000000000000000000000010110",
"000000000000000000000000000000000011111000",
"000111000000000000000000000000000000000010",
"000101100000000000000000000000000000110000",
"000100000000000000000000000000000000111000",
"000000000000000000000000000000001100000000",
"000101100000000000000000000000000000101001",
"010000000000000000000000000111100000110011",
"000000000000000000000000000000000001111100",
"000100000000000000000000000000000010101110",
"000111000000000000000000000000000000011011",
"000100000000000000000000000000001011111000",
"000000000000000000000000000000010100000000",
"000101100000000000000000000000000000101001",
"000100000000000000000000000000000000111000",
"000000000000000000000000000000110000000000",
"000111000000000000000000000000000000111100",
"000101100000000000000000000000000000101110",
"000100000000000000000000000000001000111000",
"000100000000000000000000000000000100000101",
"000101100000000000000000000000000000111100",
"000100000000000000000000000000000000111000",
"000000000000000000000000000000011100000000",
"101111111111111111111111111111111111111111",
"000101100000000000000000000000000000101110",
"000100000000000000000000000000001001111000",
"000100000000000000000000000000000101000101",
"000101100000000000000000000000000000010100",
"000100000000000000000000000000001011111000",
"000000000000000000000000000000100000000000",
"000101100000000000000000000000000000010101",
"000100000000000000000000000000000000111000",
"000000000000000000000000000000100100000000",
"000100000000000000000000000000000100111100",
"000101100000000000000000000000000000101110",
"000000000000000000000000000000100000000000",
"000101100000000000000000000000000000010010",
"101111111111111111111111111111111111111111",
"000100000000000000000000000000001010111000",
"000100000000000000000000000000000110000101",
"000101100000000000000000000000000000010100",
"000100000000000000000000000000000000111000",
"000000000000000000000000000000010100000000",
"000101100000000000000000000000000000101001",
"101111111111111111111111111111111111111111",
"000100000000000000000000000000000101101001",
"000111000000000000000000000000000000111000",
"000000000000000000000000000000000000000010",
"000101100000000000000000000000000000110000",
"001000000000000000000000000000010011110011",
"000100000000000000000000000000000100111100",
"000100000000000000000000000000000010101110",
"000111000000000000000000000000000000010101",
"000100000000000000000000000000000000111000",
"000000000000000000000000000000110000000000",
"000101100000000000000000000000000000101001",
"000100000000000000000000000000000000111000",
"000000000000000000000000000000000100000000",
"000111000000000000000000000000000000111100",
"000101100000000000000000000000000000101110",
"000000000000000000000000000000101000000000",
"000101100000000000000000000000000000010100",
"101111111111111111111111111111111111111111",
"000000000000000000000000000000110100000000",
"000101100000000000000000000000000000101001",
"000111000000000000000000000000000000010010",
"000000000000000000000000001110000101110010",
"000100000000000000000000000000000101111100",
"000100000000000000000000000000000100101110",
"000111000000000000000000000000000000010001",
"000100000000000000000000000000000000111000",
"000000000000000000000000000000101000000000",
"000101100000000000000000000000000000101001",
"000000000000000000000000000000000000011011",
"000000000000000000000000000000000000010101",
"000111000000000000000000000000000000011100",
"000100000000000000000000000000000010111000",
"000100000000000000000000000000000010000000",
"000101100000000000000000000000000000010100",
"000100000000000000000000000000000000111000",
"000000000000000000000000000000101100000000",
"000101100000000000000000000000000000010010",
"000100000000000000000000000000000100111000",
"000100000000000000000000000000000100000000",
"000101100000000000000000000000000000111100",
"000100000000000000000000000000000010101110",
"000100000000000000000000000000000000111000",
"000000000000000000000000000000010000000000",
"000101100000000000000000000000000000010010",
"000100000000000000000000000000000001111000",
"000100000000000000000000000000000001000000",
"000101100000000000000000000000000000111000",
"000000000000000000000000001001011111110011",
"000101100000000000000000000000000000000000",
"000101100000000000000000000000000000111100",
"000100000000000000000000000000000010101110",
"000100000000000000000000000000000000111000",
"000000000000000000000000000000100000000000",
"000101100000000000000000000000000000010010",
"000000000000000000000000000000010000000000",
"000101100000000000000000000000000000101001",
"101111111111111111111111111111111111111111",
"101111111111111111111111111111111111111111",
"000000000000000000000000000000100000000000",
"000101100000000000000000000000000000101001",
"000111000000000000000000000000000000010101",
"000111000000000000000000000000000000111000",
"000111000000000000000000000000000000000000",
"000101100000000000000000000000000000111100",
"000100000000000000000000000000000010101110",
"000100000000000000000000000000000000111000",
"000000000000000000000000000000100100000000",
"000101100000000000000000000000000000010010",
"000000000000000000000000000000100100000000",
"000101100000000000000000000000000000101001",
"101111111111111111111111111111111111111111",
"101111111111111111111111111111111111111111",
"000100000000000000000000000000000101111000",
"000111000000000000000000000000000000000000",
"000101100000000000000000000000000000111100",
"000100000000000000000000000000000000111000",
"000000000000000000000000000000011100000000",
"000101100000000000000000000000000000101001",
"000100000000000000000000000000000010101110",
"000100000000000000000000000000000101111000",
"000111000000000000000000000000000000000000",
"000101100000000000000000000000000000111100",
"000100000000000000000000000000000000111000",
"000000000000000000000000000000010100000000",
"000101100000000000000000000000000000010100",
"000000000000000000000000000000011000000000",
"000101100000000000000000000000000000101001",
"101111111111111111111111111111111111111111",
"101111111111111111111111111111111111111111",
"000100000000000000000000000000000100101001",
"000111000000000000000000000000000000111000",
"000000000000000000000000000000000001000000",
"000101100000000000000000000000000000010101",
"000111000000000000000000000000000000111000",
"000101100000000000000000000000000000000010",
"000101100000000000000000000000000000110000",
"001000000000000000000000000000010011110011",
"000100000000000000000000000000000000111000",
"000000000000000000000000000000011100000000",
"000101100000000000000000000000000000101110",
"000100000000000000000000000000000000111000",
"000000000000000000000000000000011000000000",
"000101100000000000000000000000000000010010",
"000000000000000000000000000000110100000000",
"000101100000000000000000000000000000101001",
"101111111111111111111111111111111111111111",
"101111111111111111111111111111111111111111",
"000111000000000000000000000000000000111000",
"101111111111111111111111111111111111111111",
"000000000000000000000000000000000001000011",
"000101100000000000000000000000000000110000",
"001000000000000000000000001000101110110011",
"101111111111111111111111111111111111111111",
"000100000000000000000000000000000101111100",
"000100000000000000000000000000000010101110",
"000100000000000000000000000000000000111000",
"000000000000000000000000000000110000000000",
"000101100000000000000000000000000000101001",
"101111111111111111111111111111111111111111",
"101111111111111111111111111111111111111111",
"000111000000000000000000000000000000111000",
"000000000000000000000000000000000001000011",
"000101100000000000000000000000000000110000",
"001000000000000000000000001000110001110011",
"001100000000000000000000000000000000111000",
"001000000000000000000000000000100000000000",
"001101100000000000000000000000000000010010",
"000100000000000000000000000000001100111000",
"000000000000000000000000000000000000000010",
"000101100000000000000000000000000000110000",
"001000000000000000000000001101001110110011",
"000100000000000000000000000000000000111000",
"000000000000000000000000000000100000000000",
"000101100000000000000000000000000000010010",
"000100000000000000000000000000000010101001",
"000100000000000000000000000000000000111000",
"000000000000000000000000000001000100000000",
"000111000000000000000000000000000000111100",
"000101100000000000000000000000000000101110",
"000000000000000000000000000000100100000000",
"000101100000000000000000000000000000101001",
"101111111111111111111111111111111111111111",
"000100000000000000000000000000000000111000",
"000000000000000000000000000001000000000000",
"000111000000000000000000000000000000111100",
"000101100000000000000000000000000000101110",
"000000000000000000000000000000111100000000",
"000101100000000000000000000000000000010010",
"101111111111111111111111111111111111111111",
"000000000000000000000000000000011100000000",
"000101100000000000000000000000000000101001",
"101111111111111111111111111111111111111111",
"000000000000000000000000001011001010110011",
"000111000000000000000000000000000000111100",
"000100000000000000000000000000000010101110",
"000100000000000000000000000000001011010101",
"000100000000000000000000000000000000111000",
"000000000000000000000000000001000100000000",
"000101100000000000000000000000000000010010",
"000000000000000000000000000000101100000000",
"000101100000000000000000000000000000101001",
"000100000000000000000000000000000000111000",
"000000000000000000000000000001000100000000",
"000101100000000000000000000000000000101001",
"000111000000000000000000000000000000010100",
"000111000000000000000000000000000000111000",
"000111000000000000000000000000000000000000",
"000101100000000000000000000000000000111100",
"000100000000000000000000000000000010101110",
"000100000000000000000000000000000000111000",
"000000000000000000000000000001000000000000",
"000101100000000000000000000000000000010010",
"000000000000000000000000000000101000000000",
"000101100000000000000000000000000000101001",
"101111111111111111111111111111111111111111",
"000000000000000000000000000001000000000000",
"000101100000000000000000000000000000101001",
"000111000000000000000000000000000000011100",
"101111111111111111111111111111111111111111",
"000100000000000000000000000000000100111000",
"000111000000000000000000000000000000000000",
"000101100000000000000000000000000000010101",
"000100000000000000000000000000000000111000",
"000000000000000000000000000000111100000000",
"000101100000000000000000000000000000101001",
"000100000000000000000000000000000101111100",
"000100000000000000000000000000000100111000",
"000111000000000000000000000000000000000000",
"000101100000000000000000000000000000010101",
"000100000000000000000000000000000000111000",
"000000000000000000000000000000110100000000",
"000101100000000000000000000000000000010100",
"000000000000000000000000000000111000000000",
"000101100000000000000000000000000000101001",
"000100000000000000000000000000000010101110",
"000100000000000000000000000000000101111100",
"000100000000000000000000000000000100101001",
"000111000000000000000000000000000000111000",
"000000000000000000000000000000000001000000",
"000101100000000000000000000000000000010101",
"000111000000000000000000000000000000111000",
"000101100000000000000000000000000000000010",
"000101100000000000000000000000000000110000",
"001000000000000000000000001000101110110011",
"000100000000000000000000000000000000111000",
"000000000000000000000000000000111100000000",
"000101100000000000000000000000000000101110",
"000100000000000000000000000000001100111000",
"000000000000000000000000000000000001000010",
"000101100000000000000000000000000000110000",
"000100000000000000000000000000000000111000",
"001000000000000000000000001100011101110011",
"000000000000000000000000000000111000000000",
"000100000000000000000000000000000101111100",
"000101100000000000000000000000000000101110",
"000000000000000000000000000000000010111000",
"000100000000000000000000000000001100000010",
"000101100000000000000000000000000000110000",
"000100000000000000000000000000000000111000",
"000000000000000000000000000000110000000000",
"000101100000000000000000000000000000101001",
"000000000000000000000000000000111100000000",
"101111111111111111111111111111111111111111",
"000101100000000000000000000000000000101001",
"000000000000000000000000000001000000000000",
"000111000000000000000000000000000000010010",
"000101100000000000000000000000000000101001",
"000000000000000000000000000001000100000000",
"000111000000000000000000000000000000010111",
"000101100000000000000000000000000000101001",
"010000000000000000000000001010010111110011",
"000111000000000000000000000000000000010110",
"101111111111111111111111111111111111111111",
"000111000000000000000000000000000000010101",
"000100000000000000000000000000000000111000",
"000000000000000000000000000001001000000000",
"000100000000000000000000000000000111111100",
"000101100000000000000000000000000000101110",
"000000000000000000000000000001001100000000",
"101111111111111111111111111111111111111111",
"000100000000000000000000000000000110111100",
"000101100000000000000000000000000000101110",
"000000000000000000000000000001010000000000",
"101111111111111111111111111111111111111111",
"000100000000000000000000000000000101111100",
"000101100000000000000000000000000000101110",
"000000000000000000000000000001010000000000",
"000101100000000000000000000000000000101001",
"101111111111111111111111111111111111111111",
"000000000000000000000000000000000100000000",
"000111000000000000000000000000000000100001",
"000100000000000000000000000000000110100001",
"000000000000000000000000001110000101110010",
"000101000000000000000000000000000000111100",
"000101000000000000000000000000000000010001",
"000101100000000000000000000000000000101110",
"000100000000000000000000000000000000111000",
"000000000000000000000000000001001000000000",
"000101100000000000000000000000000000101001",
"000000000000000000000000000001001100000000",
"101111111111111111111111111111111111111111",
"000101100000000000000000000000000000101001",
"000000000000000000000000000000000000011011",
"000111000000000000000000000000000000010111",
"000111000000000000000000000000000000010110",
"000100000000000000000000000000000000111000",
"000000000000000000000000000001010000000000",
"000101100000000000000000000000000000101001",
"000100000000000000000000000000000010111000",
"000011111111111111111111111111111111000000",
"000101100000000000000000000000000000010010",
"000000000000000000000000000000000000111000",
"000101100000000000000000000000000000000010",
"000101100000000000000000000000000000110000",
"000100000000000000000000000000000001110110",
"000100000000000000000000000000000111100110",
"000100000000000000000000000000000111111000",
"000000000000000000000000000000000100000000",
"000101100000000000000000000000000000010111",
"000100000000000000000000000000000110111000",
"000000000000000000000000000000000100000000",
"000101100000000000000000000000000000010110",
"010000000000000000000000001011100101110011",
"000111000000000000000000000000000000111000",
"000000000000000000000000000000000100000000",
"000101100000000000000000000000000000010101",
"000000000000000000000000001010011001110011",
"101111111111111111111111111111111111111111",
"000100000000000000000000000000000000111000",
"000000000000000000000000000001000100000000",
"000100000000000000000000000000000000111000",
"000000000000000000000000000000110000000000",
"000101100000000000000000000000000000101001",
"101111111111111111111111111111111111111111",
"000100000000000000000000000000001011010101",
"000111000000000000000000000000000000010100",
"000100000000000000000000000000000000111000",
"000000000000000000000000000001000000000000",
"000101100000000000000000000000000000101001",
"101111111111111111111111111111111111111111",
"000100000000000000000000000000000101111000",
"000111000000000000000000000000000000000000",
"000101100000000000000000000000000000010111",
"000100000000000000000000000000000000111000",
"000000000000000000000000000001000100000000",
"000101100000000000000000000000000000101001",
"101111111111111111111111111111111111111111",
"000100000000000000000000000000000101111000",
"000111000000000000000000000000000000000000",
"000101100000000000000000000000000000100001",
"000100000000000000000000000000000111100001",
"101111111111111111111111111111111111111111",
"000101000000000000000000000000000000111000",
"000101000000000000000000000000000000000000",
"000101100000000000000000000000000000010110",
"000100000000000000000000000000000000111000",
"000000000000000000000000000000111100000000",
"000101100000000000000000000000000000101001",
"101111111111111111111111111111111111111111",
"000100000000000000000000000000000101111000",
"000111000000000000000000000000000000000000",
"000101100000000000000000000000000000010111",
"000000000000000000000000000000000100000000",
"000101100000000000000000000000000000010101",
"101111111111111111111111111111111111111111",
"000100000000000000000000000000000100111000",
"000011111111111111111111111111111111000000",
"000101100000000000000000000000000000010100",
"000101100000000000000000000000000000111000",
"000000000000000000000000000000000000000010",
"000101100000000000000000000000000000110000",
"010000000000000000000000001100100011110011",
"101111111111111111111111111111111111111111",
"000100000000000000000000000000000110110110",
"000100000000000000000000000000000111100110",
"000000000000000000000000001010011001110011",
"101111111111111111111111111111111111111111",
"000100000000000000000000000000000000111000",
"000000000000000000000000000001000100000000",
"000100000000000000000000000000000010101001",
"000100000000000000000000000000000000111000",
"000000000000000000000000000000100100000000",
"000101100000000000000000000000000000101001",
"000100000000000000000000000000001011010110",
"000111000000000000000000000000000000010100",
"000111000000000000000000000000000000010101",
"000100000000000000000000000000000000111000",
"000000000000000000000000000000110000000000",
"000101100000000000000000000000000000101001",
"000100000000000000000000000000000101011000",
"000100000000000000000000000000000100010111",
"000111000000000000000000000000000000011001",
"000100000000000000000000000000000111100001",
"000100000000000000000000000000000111111000",
"000000000000000000000000000000000100000000",
"000101100000000000000000000000000000010111",
"000101000000000000000000000000000000110110",
"000100000000000000000000000000001000100110",
"000100000000000000000000000000001001111000",
"000011111111111111111111111111111111000000",
"000101100000000000000000000000000000011001",
"000100000000000000000000000000001011111000",
"000101100000000000000000000000000000000010",
"000101100000000000000000000000000000110000",
"010000000000000000000000001101011011110011",
"000100000000000000000000000000001000111000",
"000000000000000000000000000000000100000000",
"000101100000000000000000000000000000011000",
"000100000000000000000000000000000000111000",
"000000000000000000000000000000101100000000",
"000101100000000000000000000000000000101001",
"101111111111111111111111111111111111111111",
"101111111111111111111111111111111111111111",
"000111000000000000000000000000000000010111",
"000111000000000000000000000000000000111000",
"000100000000000000000000000000000101000000",
"000101100000000000000000000000000000010101",
"000100000000000000000000000000000000111000",
"000000000000000000000000000000110100000000",
"000100000000000000000000000000000110111000",
"000101100000000000000000000000000000101001",
"000000000000000000000000000000000001000000",
"000101100000000000000000000000000000010110",
"000111000000000000000000000000000000111000",
"000101100000000000000000000000000000000010",
"000101100000000000000000000000000000110000",
"010000000000000000000000001101010101110011",
"000100000000000000000000000000000111111000",
"000100000000000000000000000000000100000000",
"000101100000000000000000000000000000010100",
"000000000000000000000000001000110000110011",
"101111111111111111111111111111111111111111",
"000100000000000000000000000000000000111000",
"000000000000000000000000000000100000000000",
"000100000000000000000000000000000001111000",
"000000000000000000000000000000000000000010",
"000101100000000000000000000000000000110000",
"001110000000000000000000000000000000110011",
"101111111111111111111111111111111111111111",
"101111111111111111111111111111111111111111",
"001000000000000000000000000000000000010001",
"000100000000000000000000000000000000111000",
"000000000000000000000000000000000100000000",
"000101100000000000000000000000000000101001",
"000000000000000000000000000000000000010110",
"000000000000000000000000000000000000010100",
"000111000000000000000000000000000000010101",
"000100000000000000000000000000000001111000",
"000000000000000000000000000000000001000001",
"000101100000000000000000000000000000111000",
"000000000000000000000000000000000000001000",
"000100000000000000000000000000000101111000",
"000101100000000000000000000000000000000001",
"000101100000000000000000000000000000010111",
"000100000000000000000000000000000101000000",
"000101100000000000000000000000000000010101",
"101111111111111111111111111111111111111111",
"000100000000000000000000000000000001000111",
"000101100000000000000000000000000000010001",
"000100000000000000000000000000000110111000",
"000101100000000000000000000000000000000010",
"000101100000000000000000000000000000110000",
"010000000000000000000000001110010010110011",
"000100000000000000000000000000000100111000",
"000100000000000000000000000000000111000000",
"000101100000000000000000000000000000010100",
"000110000000000000000000000000000000110011",
"101111111111111111111111111111111111111111",
"101111111111111111111111111111111111111111",
"000100000000000000000000000000000100010001");

end tta_core_imem_image;

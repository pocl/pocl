package tta_core_params is
end tta_core_params;

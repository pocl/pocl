package ffaccel_params is
  constant fu_DATA_LSU_addrw_g : integer := 12;
  constant fu_PARAM_LSU_addrw_g : integer := 32;
  constant fu_SP_LSU_addrw_g : integer := 10;
end ffaccel_params;

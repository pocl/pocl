package tta_core_toplevel_params is
end tta_core_toplevel_params;

package ffaccel_imem_mau is
   -- created by generatebits
   constant IMEMMAUWIDTH : positive := 43;
end ffaccel_imem_mau;
